BZh91AY&SYu��I _�Px�w��߰?���Px=;��ց��T�h��2z	���� OH?T�5=&F�0#A��ɑ��hdb��&��F��jm50��4  bb=M4�ɓF�� �0F`H�4 F)?"�=#j4�@��H|�h�J�BC:�>=T[F��؁�t�ҀX1�af����0H����}$��Ba�l�]���IR)�/�A����L��&���2*�G=���e>���h���n���l�Ci:���"m�E�&)�u��,���tr�ʲa�����]�D_���g�wt�+5�)pВ�
'=N�0Q����h�Ï(ʄ%q�`Q��h
 x�8��atD��|͙a�=�u�'�c�t�j���EJ���Ҁ{�'��S�YH˰������xh��;$�/*6�<WE���.N�ي�[!������Ő^���`t�*qz]5�i����M�r�o<���>ǯ��DF<L樓�'l��gE
�m3#n�4��I3��n`y@t%`�yR�J1ߐ?���7޻P��eʧG�7I�\mOMϰ�T3��P0��-��˺.��o��a=̤;A��o�7����:�)V�}�ʸ�r%�2�H�D`�����p�p4��0��Ic��
/���@�~�TXNťp�(��rg�4�_j99A�3�U�.q�9W��s�M�� ����Ⱥ9�a��TM���TR��3q�$�?��S"`���BDZ餏܎=8�D�Jl�hH��K6`�O|�΂�S-Jc�F���x�)����F���kQ,r.�M���d�e�1�fd���D��"�(H:�V$�